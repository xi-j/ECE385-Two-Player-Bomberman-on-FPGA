// Bomberman.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Bomberman (
		output wire [7:0]  audio_back_vol_export,     //     audio_back_vol.export
		output wire        audio_bomb_active_export,  //  audio_bomb_active.export
		output wire [2:0]  audio_bomb_vol_export,     //     audio_bomb_vol.export
		output wire        audio_init_export,         //         audio_init.export
		input  wire        audio_init_f_export,       //       audio_init_f.export
		output wire [2:0]  audio_select_export,       //       audio_select.export
		input  wire        boot_up_export,            //            boot_up.export
		input  wire        clk_clk,                   //                clk.clk
		output wire [8:0]  export_data_new_signal,    //        export_data.new_signal
		output wire [31:0] export_data_new_signal_1,  //                   .new_signal_1
		output wire [63:0] export_data_new_signal_2,  //                   .new_signal_2
		input  wire        export_data_new_signal_3,  //                   .new_signal_3
		output wire        export_data_new_signal_4,  //                   .new_signal_4
		output wire [7:0]  led_wire_export,           //           led_wire.export
		output wire [1:0]  otg_hpi_address_export,    //    otg_hpi_address.export
		output wire        otg_hpi_cs_export,         //         otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,      //       otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,     //                   .out_port
		output wire        otg_hpi_r_export,          //          otg_hpi_r.export
		output wire        otg_hpi_reset_export,      //      otg_hpi_reset.export
		output wire        otg_hpi_w_export,          //          otg_hpi_w.export
		output wire [3:0]  player1score0_wire_export, // player1score0_wire.export
		output wire [3:0]  player1score1_wire_export, // player1score1_wire.export
		output wire [3:0]  player2score0_wire_export, // player2score0_wire.export
		output wire [3:0]  player2score1_wire_export, // player2score1_wire.export
		input  wire        reset_reset_n,             //              reset.reset_n
		output wire        sdram_pll_clk,             //          sdram_pll.clk
		output wire [12:0] sdram_wire_addr,           //         sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,             //                   .ba
		output wire        sdram_wire_cas_n,          //                   .cas_n
		output wire        sdram_wire_cke,            //                   .cke
		output wire        sdram_wire_cs_n,           //                   .cs_n
		inout  wire [31:0] sdram_wire_dq,             //                   .dq
		output wire [3:0]  sdram_wire_dqm,            //                   .dqm
		output wire        sdram_wire_ras_n,          //                   .ras_n
		output wire        sdram_wire_we_n,           //                   .we_n
		output wire [3:0]  timescreen0_wire_export,   //   timescreen0_wire.export
		output wire [3:0]  timescreen1_wire_export,   //   timescreen1_wire.export
		output wire [3:0]  timescreen2_wire_export    //   timescreen2_wire.export
	);

	wire         sdram_pll_audio_pll_c0_clk;                                  // sdram_pll_audio_pll:c0 -> [mm_interconnect_0:sdram_pll_audio_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                        // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [27:0] nios2_qsys_0_data_master_address;                            // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                         // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                               // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                              // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                          // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [27:0] nios2_qsys_0_instruction_master_address;                     // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                        // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;     // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;  // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_audio_pll_pll_slave_readdata;    // sdram_pll_audio_pll:readdata -> mm_interconnect_0:sdram_pll_audio_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_audio_pll_pll_slave_address;     // mm_interconnect_0:sdram_pll_audio_pll_pll_slave_address -> sdram_pll_audio_pll:address
	wire         mm_interconnect_0_sdram_pll_audio_pll_pll_slave_read;        // mm_interconnect_0:sdram_pll_audio_pll_pll_slave_read -> sdram_pll_audio_pll:read
	wire         mm_interconnect_0_sdram_pll_audio_pll_pll_slave_write;       // mm_interconnect_0:sdram_pll_audio_pll_pll_slave_write -> sdram_pll_audio_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_audio_pll_pll_slave_writedata;   // mm_interconnect_0:sdram_pll_audio_pll_pll_slave_writedata -> sdram_pll_audio_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_avalon_blitter_0_s1_chipselect;            // mm_interconnect_0:avalon_blitter_0_s1_chipselect -> avalon_blitter_0:AVL_CS
	wire  [31:0] mm_interconnect_0_avalon_blitter_0_s1_readdata;              // avalon_blitter_0:AVL_READDATA -> mm_interconnect_0:avalon_blitter_0_s1_readdata
	wire   [4:0] mm_interconnect_0_avalon_blitter_0_s1_address;               // mm_interconnect_0:avalon_blitter_0_s1_address -> avalon_blitter_0:AVL_ADDR
	wire         mm_interconnect_0_avalon_blitter_0_s1_read;                  // mm_interconnect_0:avalon_blitter_0_s1_read -> avalon_blitter_0:AVL_READ
	wire   [3:0] mm_interconnect_0_avalon_blitter_0_s1_byteenable;            // mm_interconnect_0:avalon_blitter_0_s1_byteenable -> avalon_blitter_0:AVL_BYTE_EN
	wire         mm_interconnect_0_avalon_blitter_0_s1_write;                 // mm_interconnect_0:avalon_blitter_0_s1_write -> avalon_blitter_0:AVL_WRITE
	wire  [31:0] mm_interconnect_0_avalon_blitter_0_s1_writedata;             // mm_interconnect_0:avalon_blitter_0_s1_writedata -> avalon_blitter_0:AVL_WRITEDATA
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;               // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                 // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                  // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                    // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_audio_init_s1_chipselect;                  // mm_interconnect_0:audio_INIT_s1_chipselect -> audio_INIT:chipselect
	wire  [31:0] mm_interconnect_0_audio_init_s1_readdata;                    // audio_INIT:readdata -> mm_interconnect_0:audio_INIT_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_init_s1_address;                     // mm_interconnect_0:audio_INIT_s1_address -> audio_INIT:address
	wire         mm_interconnect_0_audio_init_s1_write;                       // mm_interconnect_0:audio_INIT_s1_write -> audio_INIT:write_n
	wire  [31:0] mm_interconnect_0_audio_init_s1_writedata;                   // mm_interconnect_0:audio_INIT_s1_writedata -> audio_INIT:writedata
	wire  [31:0] mm_interconnect_0_audio_init_f_s1_readdata;                  // audio_INIT_F:readdata -> mm_interconnect_0:audio_INIT_F_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_init_f_s1_address;                   // mm_interconnect_0:audio_INIT_F_s1_address -> audio_INIT_F:address
	wire         mm_interconnect_0_audio_back_vol_s1_chipselect;              // mm_interconnect_0:audio_back_vol_s1_chipselect -> audio_back_vol:chipselect
	wire  [31:0] mm_interconnect_0_audio_back_vol_s1_readdata;                // audio_back_vol:readdata -> mm_interconnect_0:audio_back_vol_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_back_vol_s1_address;                 // mm_interconnect_0:audio_back_vol_s1_address -> audio_back_vol:address
	wire         mm_interconnect_0_audio_back_vol_s1_write;                   // mm_interconnect_0:audio_back_vol_s1_write -> audio_back_vol:write_n
	wire  [31:0] mm_interconnect_0_audio_back_vol_s1_writedata;               // mm_interconnect_0:audio_back_vol_s1_writedata -> audio_back_vol:writedata
	wire         mm_interconnect_0_audio_bomb_vol_s1_chipselect;              // mm_interconnect_0:audio_bomb_vol_s1_chipselect -> audio_bomb_vol:chipselect
	wire  [31:0] mm_interconnect_0_audio_bomb_vol_s1_readdata;                // audio_bomb_vol:readdata -> mm_interconnect_0:audio_bomb_vol_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_bomb_vol_s1_address;                 // mm_interconnect_0:audio_bomb_vol_s1_address -> audio_bomb_vol:address
	wire         mm_interconnect_0_audio_bomb_vol_s1_write;                   // mm_interconnect_0:audio_bomb_vol_s1_write -> audio_bomb_vol:write_n
	wire  [31:0] mm_interconnect_0_audio_bomb_vol_s1_writedata;               // mm_interconnect_0:audio_bomb_vol_s1_writedata -> audio_bomb_vol:writedata
	wire         mm_interconnect_0_audio_bomb_active_s1_chipselect;           // mm_interconnect_0:audio_bomb_active_s1_chipselect -> audio_bomb_active:chipselect
	wire  [31:0] mm_interconnect_0_audio_bomb_active_s1_readdata;             // audio_bomb_active:readdata -> mm_interconnect_0:audio_bomb_active_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_bomb_active_s1_address;              // mm_interconnect_0:audio_bomb_active_s1_address -> audio_bomb_active:address
	wire         mm_interconnect_0_audio_bomb_active_s1_write;                // mm_interconnect_0:audio_bomb_active_s1_write -> audio_bomb_active:write_n
	wire  [31:0] mm_interconnect_0_audio_bomb_active_s1_writedata;            // mm_interconnect_0:audio_bomb_active_s1_writedata -> audio_bomb_active:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_player2score0_s1_chipselect;               // mm_interconnect_0:player2Score0_s1_chipselect -> player2Score0:chipselect
	wire  [31:0] mm_interconnect_0_player2score0_s1_readdata;                 // player2Score0:readdata -> mm_interconnect_0:player2Score0_s1_readdata
	wire   [1:0] mm_interconnect_0_player2score0_s1_address;                  // mm_interconnect_0:player2Score0_s1_address -> player2Score0:address
	wire         mm_interconnect_0_player2score0_s1_write;                    // mm_interconnect_0:player2Score0_s1_write -> player2Score0:write_n
	wire  [31:0] mm_interconnect_0_player2score0_s1_writedata;                // mm_interconnect_0:player2Score0_s1_writedata -> player2Score0:writedata
	wire         mm_interconnect_0_player2score1_s1_chipselect;               // mm_interconnect_0:player2Score1_s1_chipselect -> player2Score1:chipselect
	wire  [31:0] mm_interconnect_0_player2score1_s1_readdata;                 // player2Score1:readdata -> mm_interconnect_0:player2Score1_s1_readdata
	wire   [1:0] mm_interconnect_0_player2score1_s1_address;                  // mm_interconnect_0:player2Score1_s1_address -> player2Score1:address
	wire         mm_interconnect_0_player2score1_s1_write;                    // mm_interconnect_0:player2Score1_s1_write -> player2Score1:write_n
	wire  [31:0] mm_interconnect_0_player2score1_s1_writedata;                // mm_interconnect_0:player2Score1_s1_writedata -> player2Score1:writedata
	wire         mm_interconnect_0_player1score0_s1_chipselect;               // mm_interconnect_0:player1Score0_s1_chipselect -> player1Score0:chipselect
	wire  [31:0] mm_interconnect_0_player1score0_s1_readdata;                 // player1Score0:readdata -> mm_interconnect_0:player1Score0_s1_readdata
	wire   [1:0] mm_interconnect_0_player1score0_s1_address;                  // mm_interconnect_0:player1Score0_s1_address -> player1Score0:address
	wire         mm_interconnect_0_player1score0_s1_write;                    // mm_interconnect_0:player1Score0_s1_write -> player1Score0:write_n
	wire  [31:0] mm_interconnect_0_player1score0_s1_writedata;                // mm_interconnect_0:player1Score0_s1_writedata -> player1Score0:writedata
	wire         mm_interconnect_0_player1score1_s1_chipselect;               // mm_interconnect_0:player1Score1_s1_chipselect -> player1Score1:chipselect
	wire  [31:0] mm_interconnect_0_player1score1_s1_readdata;                 // player1Score1:readdata -> mm_interconnect_0:player1Score1_s1_readdata
	wire   [1:0] mm_interconnect_0_player1score1_s1_address;                  // mm_interconnect_0:player1Score1_s1_address -> player1Score1:address
	wire         mm_interconnect_0_player1score1_s1_write;                    // mm_interconnect_0:player1Score1_s1_write -> player1Score1:write_n
	wire  [31:0] mm_interconnect_0_player1score1_s1_writedata;                // mm_interconnect_0:player1Score1_s1_writedata -> player1Score1:writedata
	wire         mm_interconnect_0_timescreen1_s1_chipselect;                 // mm_interconnect_0:timeScreen1_s1_chipselect -> timeScreen1:chipselect
	wire  [31:0] mm_interconnect_0_timescreen1_s1_readdata;                   // timeScreen1:readdata -> mm_interconnect_0:timeScreen1_s1_readdata
	wire   [1:0] mm_interconnect_0_timescreen1_s1_address;                    // mm_interconnect_0:timeScreen1_s1_address -> timeScreen1:address
	wire         mm_interconnect_0_timescreen1_s1_write;                      // mm_interconnect_0:timeScreen1_s1_write -> timeScreen1:write_n
	wire  [31:0] mm_interconnect_0_timescreen1_s1_writedata;                  // mm_interconnect_0:timeScreen1_s1_writedata -> timeScreen1:writedata
	wire         mm_interconnect_0_timescreen2_s1_chipselect;                 // mm_interconnect_0:timeScreen2_s1_chipselect -> timeScreen2:chipselect
	wire  [31:0] mm_interconnect_0_timescreen2_s1_readdata;                   // timeScreen2:readdata -> mm_interconnect_0:timeScreen2_s1_readdata
	wire   [1:0] mm_interconnect_0_timescreen2_s1_address;                    // mm_interconnect_0:timeScreen2_s1_address -> timeScreen2:address
	wire         mm_interconnect_0_timescreen2_s1_write;                      // mm_interconnect_0:timeScreen2_s1_write -> timeScreen2:write_n
	wire  [31:0] mm_interconnect_0_timescreen2_s1_writedata;                  // mm_interconnect_0:timeScreen2_s1_writedata -> timeScreen2:writedata
	wire         mm_interconnect_0_timescreen0_s1_chipselect;                 // mm_interconnect_0:timeScreen0_s1_chipselect -> timeScreen0:chipselect
	wire  [31:0] mm_interconnect_0_timescreen0_s1_readdata;                   // timeScreen0:readdata -> mm_interconnect_0:timeScreen0_s1_readdata
	wire   [1:0] mm_interconnect_0_timescreen0_s1_address;                    // mm_interconnect_0:timeScreen0_s1_address -> timeScreen0:address
	wire         mm_interconnect_0_timescreen0_s1_write;                      // mm_interconnect_0:timeScreen0_s1_write -> timeScreen0:write_n
	wire  [31:0] mm_interconnect_0_timescreen0_s1_writedata;                  // mm_interconnect_0:timeScreen0_s1_writedata -> timeScreen0:writedata
	wire         mm_interconnect_0_audio_select_s1_chipselect;                // mm_interconnect_0:audio_select_s1_chipselect -> audio_select:chipselect
	wire  [31:0] mm_interconnect_0_audio_select_s1_readdata;                  // audio_select:readdata -> mm_interconnect_0:audio_select_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_select_s1_address;                   // mm_interconnect_0:audio_select_s1_address -> audio_select:address
	wire         mm_interconnect_0_audio_select_s1_write;                     // mm_interconnect_0:audio_select_s1_write -> audio_select:write_n
	wire  [31:0] mm_interconnect_0_audio_select_s1_writedata;                 // mm_interconnect_0:audio_select_s1_writedata -> audio_select:writedata
	wire  [31:0] mm_interconnect_0_boot_up_s1_readdata;                       // Boot_Up:readdata -> mm_interconnect_0:Boot_Up_s1_readdata
	wire   [1:0] mm_interconnect_0_boot_up_s1_address;                        // mm_interconnect_0:Boot_Up_s1_address -> Boot_Up:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Boot_Up:reset_n, LEDs:reset_n, audio_INIT:reset_n, audio_INIT_F:reset_n, audio_back_vol:reset_n, audio_bomb_active:reset_n, audio_bomb_vol:reset_n, audio_select:reset_n, mm_interconnect_0:sdram_pll_audio_pll_inclk_interface_reset_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, player1Score0:reset_n, player1Score1:reset_n, player2Score0:reset_n, player2Score1:reset_n, sdram_pll_audio_pll:reset, timeScreen0:reset_n, timeScreen1:reset_n, timeScreen2:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [avalon_blitter_0:Hard_RESET, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                      // nios2_qsys_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	Bomberman_Boot_Up boot_up (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_boot_up_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boot_up_s1_readdata), //                    .readdata
		.in_port  (boot_up_export)                         // external_connection.export
	);

	Bomberman_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (led_wire_export)                       // external_connection.export
	);

	Bomberman_audio_INIT audio_init (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_audio_init_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_init_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_init_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_init_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_init_s1_readdata),   //                    .readdata
		.out_port   (audio_init_export)                           // external_connection.export
	);

	Bomberman_Boot_Up audio_init_f (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_audio_init_f_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_audio_init_f_s1_readdata), //                    .readdata
		.in_port  (audio_init_f_export)                         // external_connection.export
	);

	Bomberman_LEDs audio_back_vol (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_audio_back_vol_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_back_vol_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_back_vol_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_back_vol_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_back_vol_s1_readdata),   //                    .readdata
		.out_port   (audio_back_vol_export)                           // external_connection.export
	);

	Bomberman_audio_INIT audio_bomb_active (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_audio_bomb_active_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_bomb_active_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_bomb_active_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_bomb_active_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_bomb_active_s1_readdata),   //                    .readdata
		.out_port   (audio_bomb_active_export)                           // external_connection.export
	);

	Bomberman_audio_bomb_vol audio_bomb_vol (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_audio_bomb_vol_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_bomb_vol_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_bomb_vol_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_bomb_vol_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_bomb_vol_s1_readdata),   //                    .readdata
		.out_port   (audio_bomb_vol_export)                           // external_connection.export
	);

	Bomberman_audio_bomb_vol audio_select (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_audio_select_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_select_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_select_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_select_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_select_s1_readdata),   //                    .readdata
		.out_port   (audio_select_export)                           // external_connection.export
	);

	avalon_blitter_interface avalon_blitter_0 (
		.CLOCK               (clk_clk),                                          //    clk.clk
		.AVL_ADDR            (mm_interconnect_0_avalon_blitter_0_s1_address),    //     s1.address
		.AVL_READ            (mm_interconnect_0_avalon_blitter_0_s1_read),       //       .read
		.AVL_WRITE           (mm_interconnect_0_avalon_blitter_0_s1_write),      //       .write
		.AVL_CS              (mm_interconnect_0_avalon_blitter_0_s1_chipselect), //       .chipselect
		.AVL_READDATA        (mm_interconnect_0_avalon_blitter_0_s1_readdata),   //       .readdata
		.AVL_WRITEDATA       (mm_interconnect_0_avalon_blitter_0_s1_writedata),  //       .writedata
		.AVL_BYTE_EN         (mm_interconnect_0_avalon_blitter_0_s1_byteenable), //       .byteenable
		.EXPORT_DATA         (export_data_new_signal),                           // Export.new_signal
		.EXPORT_TEST         (export_data_new_signal_1),                         //       .new_signal_1
		.Data_to_Blitter     (export_data_new_signal_2),                         //       .new_signal_2
		.Blitter_Finish_Flip (export_data_new_signal_3),                         //       .new_signal_3
		.Status_REG_Out      (export_data_new_signal_4),                         //       .new_signal_4
		.Hard_RESET          (rst_controller_001_reset_out_reset)                //  RESET.reset
	);

	Bomberman_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	Bomberman_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	Bomberman_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	Bomberman_audio_INIT otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	Bomberman_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	Bomberman_audio_INIT otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	Bomberman_audio_INIT otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	Bomberman_audio_INIT otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	Bomberman_player1Score0 player1score0 (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_player1score0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_player1score0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_player1score0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_player1score0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_player1score0_s1_readdata),   //                    .readdata
		.out_port   (player1score0_wire_export)                      // external_connection.export
	);

	Bomberman_player1Score0 player1score1 (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_player1score1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_player1score1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_player1score1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_player1score1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_player1score1_s1_readdata),   //                    .readdata
		.out_port   (player1score1_wire_export)                      // external_connection.export
	);

	Bomberman_player1Score0 player2score0 (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_player2score0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_player2score0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_player2score0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_player2score0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_player2score0_s1_readdata),   //                    .readdata
		.out_port   (player2score0_wire_export)                      // external_connection.export
	);

	Bomberman_player1Score0 player2score1 (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_player2score1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_player2score1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_player2score1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_player2score1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_player2score1_s1_readdata),   //                    .readdata
		.out_port   (player2score1_wire_export)                      // external_connection.export
	);

	Bomberman_sdram sdram (
		.clk            (sdram_pll_audio_pll_c0_clk),               //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Bomberman_sdram_pll_audio_pll sdram_pll_audio_pll (
		.clk                (clk_clk),                                                   //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                            // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_audio_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_pll_clk),                                             //                    c1.clk
		.c2                 (),                                                          //                    c2.clk
		.c3                 (),                                                          //                    c3.clk
		.scandone           (),                                                          //           (terminated)
		.scandataout        (),                                                          //           (terminated)
		.areset             (1'b0),                                                      //           (terminated)
		.locked             (),                                                          //           (terminated)
		.phasedone          (),                                                          //           (terminated)
		.phasecounterselect (4'b0000),                                                   //           (terminated)
		.phaseupdown        (1'b0),                                                      //           (terminated)
		.phasestep          (1'b0),                                                      //           (terminated)
		.scanclk            (1'b0),                                                      //           (terminated)
		.scanclkena         (1'b0),                                                      //           (terminated)
		.scandata           (1'b0),                                                      //           (terminated)
		.configupdate       (1'b0)                                                       //           (terminated)
	);

	Bomberman_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	Bomberman_player1Score0 timescreen0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_timescreen0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timescreen0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timescreen0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timescreen0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timescreen0_s1_readdata),   //                    .readdata
		.out_port   (timescreen0_wire_export)                      // external_connection.export
	);

	Bomberman_player1Score0 timescreen1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_timescreen1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timescreen1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timescreen1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timescreen1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timescreen1_s1_readdata),   //                    .readdata
		.out_port   (timescreen1_wire_export)                      // external_connection.export
	);

	Bomberman_player1Score0 timescreen2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_timescreen2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timescreen2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timescreen2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timescreen2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timescreen2_s1_readdata),   //                    .readdata
		.out_port   (timescreen2_wire_export)                      // external_connection.export
	);

	Bomberman_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	Bomberman_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                         (clk_clk),                                                     //                                                       clk_0_clk.clk
		.sdram_pll_audio_pll_c0_clk                                            (sdram_pll_audio_pll_c0_clk),                                  //                                          sdram_pll_audio_pll_c0.clk
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset                        (rst_controller_001_reset_out_reset),                          //                        nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sdram_pll_audio_pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // sdram_pll_audio_pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                               (rst_controller_002_reset_out_reset),                          //                               sdram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                                      (nios2_qsys_0_data_master_address),                            //                                        nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                                  (nios2_qsys_0_data_master_waitrequest),                        //                                                                .waitrequest
		.nios2_qsys_0_data_master_byteenable                                   (nios2_qsys_0_data_master_byteenable),                         //                                                                .byteenable
		.nios2_qsys_0_data_master_read                                         (nios2_qsys_0_data_master_read),                               //                                                                .read
		.nios2_qsys_0_data_master_readdata                                     (nios2_qsys_0_data_master_readdata),                           //                                                                .readdata
		.nios2_qsys_0_data_master_write                                        (nios2_qsys_0_data_master_write),                              //                                                                .write
		.nios2_qsys_0_data_master_writedata                                    (nios2_qsys_0_data_master_writedata),                          //                                                                .writedata
		.nios2_qsys_0_data_master_debugaccess                                  (nios2_qsys_0_data_master_debugaccess),                        //                                                                .debugaccess
		.nios2_qsys_0_instruction_master_address                               (nios2_qsys_0_instruction_master_address),                     //                                 nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                           (nios2_qsys_0_instruction_master_waitrequest),                 //                                                                .waitrequest
		.nios2_qsys_0_instruction_master_read                                  (nios2_qsys_0_instruction_master_read),                        //                                                                .read
		.nios2_qsys_0_instruction_master_readdata                              (nios2_qsys_0_instruction_master_readdata),                    //                                                                .readdata
		.audio_back_vol_s1_address                                             (mm_interconnect_0_audio_back_vol_s1_address),                 //                                               audio_back_vol_s1.address
		.audio_back_vol_s1_write                                               (mm_interconnect_0_audio_back_vol_s1_write),                   //                                                                .write
		.audio_back_vol_s1_readdata                                            (mm_interconnect_0_audio_back_vol_s1_readdata),                //                                                                .readdata
		.audio_back_vol_s1_writedata                                           (mm_interconnect_0_audio_back_vol_s1_writedata),               //                                                                .writedata
		.audio_back_vol_s1_chipselect                                          (mm_interconnect_0_audio_back_vol_s1_chipselect),              //                                                                .chipselect
		.audio_bomb_active_s1_address                                          (mm_interconnect_0_audio_bomb_active_s1_address),              //                                            audio_bomb_active_s1.address
		.audio_bomb_active_s1_write                                            (mm_interconnect_0_audio_bomb_active_s1_write),                //                                                                .write
		.audio_bomb_active_s1_readdata                                         (mm_interconnect_0_audio_bomb_active_s1_readdata),             //                                                                .readdata
		.audio_bomb_active_s1_writedata                                        (mm_interconnect_0_audio_bomb_active_s1_writedata),            //                                                                .writedata
		.audio_bomb_active_s1_chipselect                                       (mm_interconnect_0_audio_bomb_active_s1_chipselect),           //                                                                .chipselect
		.audio_bomb_vol_s1_address                                             (mm_interconnect_0_audio_bomb_vol_s1_address),                 //                                               audio_bomb_vol_s1.address
		.audio_bomb_vol_s1_write                                               (mm_interconnect_0_audio_bomb_vol_s1_write),                   //                                                                .write
		.audio_bomb_vol_s1_readdata                                            (mm_interconnect_0_audio_bomb_vol_s1_readdata),                //                                                                .readdata
		.audio_bomb_vol_s1_writedata                                           (mm_interconnect_0_audio_bomb_vol_s1_writedata),               //                                                                .writedata
		.audio_bomb_vol_s1_chipselect                                          (mm_interconnect_0_audio_bomb_vol_s1_chipselect),              //                                                                .chipselect
		.audio_INIT_s1_address                                                 (mm_interconnect_0_audio_init_s1_address),                     //                                                   audio_INIT_s1.address
		.audio_INIT_s1_write                                                   (mm_interconnect_0_audio_init_s1_write),                       //                                                                .write
		.audio_INIT_s1_readdata                                                (mm_interconnect_0_audio_init_s1_readdata),                    //                                                                .readdata
		.audio_INIT_s1_writedata                                               (mm_interconnect_0_audio_init_s1_writedata),                   //                                                                .writedata
		.audio_INIT_s1_chipselect                                              (mm_interconnect_0_audio_init_s1_chipselect),                  //                                                                .chipselect
		.audio_INIT_F_s1_address                                               (mm_interconnect_0_audio_init_f_s1_address),                   //                                                 audio_INIT_F_s1.address
		.audio_INIT_F_s1_readdata                                              (mm_interconnect_0_audio_init_f_s1_readdata),                  //                                                                .readdata
		.audio_select_s1_address                                               (mm_interconnect_0_audio_select_s1_address),                   //                                                 audio_select_s1.address
		.audio_select_s1_write                                                 (mm_interconnect_0_audio_select_s1_write),                     //                                                                .write
		.audio_select_s1_readdata                                              (mm_interconnect_0_audio_select_s1_readdata),                  //                                                                .readdata
		.audio_select_s1_writedata                                             (mm_interconnect_0_audio_select_s1_writedata),                 //                                                                .writedata
		.audio_select_s1_chipselect                                            (mm_interconnect_0_audio_select_s1_chipselect),                //                                                                .chipselect
		.avalon_blitter_0_s1_address                                           (mm_interconnect_0_avalon_blitter_0_s1_address),               //                                             avalon_blitter_0_s1.address
		.avalon_blitter_0_s1_write                                             (mm_interconnect_0_avalon_blitter_0_s1_write),                 //                                                                .write
		.avalon_blitter_0_s1_read                                              (mm_interconnect_0_avalon_blitter_0_s1_read),                  //                                                                .read
		.avalon_blitter_0_s1_readdata                                          (mm_interconnect_0_avalon_blitter_0_s1_readdata),              //                                                                .readdata
		.avalon_blitter_0_s1_writedata                                         (mm_interconnect_0_avalon_blitter_0_s1_writedata),             //                                                                .writedata
		.avalon_blitter_0_s1_byteenable                                        (mm_interconnect_0_avalon_blitter_0_s1_byteenable),            //                                                                .byteenable
		.avalon_blitter_0_s1_chipselect                                        (mm_interconnect_0_avalon_blitter_0_s1_chipselect),            //                                                                .chipselect
		.Boot_Up_s1_address                                                    (mm_interconnect_0_boot_up_s1_address),                        //                                                      Boot_Up_s1.address
		.Boot_Up_s1_readdata                                                   (mm_interconnect_0_boot_up_s1_readdata),                       //                                                                .readdata
		.jtag_uart_0_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                                   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                                .write
		.jtag_uart_0_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                                .chipselect
		.LEDs_s1_address                                                       (mm_interconnect_0_leds_s1_address),                           //                                                         LEDs_s1.address
		.LEDs_s1_write                                                         (mm_interconnect_0_leds_s1_write),                             //                                                                .write
		.LEDs_s1_readdata                                                      (mm_interconnect_0_leds_s1_readdata),                          //                                                                .readdata
		.LEDs_s1_writedata                                                     (mm_interconnect_0_leds_s1_writedata),                         //                                                                .writedata
		.LEDs_s1_chipselect                                                    (mm_interconnect_0_leds_s1_chipselect),                        //                                                                .chipselect
		.nios2_qsys_0_debug_mem_slave_address                                  (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),      //                                    nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write                                    (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),        //                                                                .write
		.nios2_qsys_0_debug_mem_slave_read                                     (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),         //                                                                .read
		.nios2_qsys_0_debug_mem_slave_readdata                                 (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),     //                                                                .readdata
		.nios2_qsys_0_debug_mem_slave_writedata                                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),    //                                                                .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable                               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),   //                                                                .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest                              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),  //                                                                .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess                              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),  //                                                                .debugaccess
		.otg_hpi_address_s1_address                                            (mm_interconnect_0_otg_hpi_address_s1_address),                //                                              otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                                              (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                                                .write
		.otg_hpi_address_s1_readdata                                           (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                                                .readdata
		.otg_hpi_address_s1_writedata                                          (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                                                .writedata
		.otg_hpi_address_s1_chipselect                                         (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                                                .chipselect
		.otg_hpi_cs_s1_address                                                 (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                                                   otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                                                   (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                                                .write
		.otg_hpi_cs_s1_readdata                                                (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                                                .readdata
		.otg_hpi_cs_s1_writedata                                               (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                                                .writedata
		.otg_hpi_cs_s1_chipselect                                              (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                                                .chipselect
		.otg_hpi_data_s1_address                                               (mm_interconnect_0_otg_hpi_data_s1_address),                   //                                                 otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                                                 (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                                                .write
		.otg_hpi_data_s1_readdata                                              (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                                                .readdata
		.otg_hpi_data_s1_writedata                                             (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                                                .writedata
		.otg_hpi_data_s1_chipselect                                            (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                                                .chipselect
		.otg_hpi_r_s1_address                                                  (mm_interconnect_0_otg_hpi_r_s1_address),                      //                                                    otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                                                    (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                                                .write
		.otg_hpi_r_s1_readdata                                                 (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                                                .readdata
		.otg_hpi_r_s1_writedata                                                (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                                                .writedata
		.otg_hpi_r_s1_chipselect                                               (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                                                .chipselect
		.otg_hpi_reset_s1_address                                              (mm_interconnect_0_otg_hpi_reset_s1_address),                  //                                                otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                                                (mm_interconnect_0_otg_hpi_reset_s1_write),                    //                                                                .write
		.otg_hpi_reset_s1_readdata                                             (mm_interconnect_0_otg_hpi_reset_s1_readdata),                 //                                                                .readdata
		.otg_hpi_reset_s1_writedata                                            (mm_interconnect_0_otg_hpi_reset_s1_writedata),                //                                                                .writedata
		.otg_hpi_reset_s1_chipselect                                           (mm_interconnect_0_otg_hpi_reset_s1_chipselect),               //                                                                .chipselect
		.otg_hpi_w_s1_address                                                  (mm_interconnect_0_otg_hpi_w_s1_address),                      //                                                    otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                                                    (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                                                .write
		.otg_hpi_w_s1_readdata                                                 (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                                                .readdata
		.otg_hpi_w_s1_writedata                                                (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                                                .writedata
		.otg_hpi_w_s1_chipselect                                               (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                                                .chipselect
		.player1Score0_s1_address                                              (mm_interconnect_0_player1score0_s1_address),                  //                                                player1Score0_s1.address
		.player1Score0_s1_write                                                (mm_interconnect_0_player1score0_s1_write),                    //                                                                .write
		.player1Score0_s1_readdata                                             (mm_interconnect_0_player1score0_s1_readdata),                 //                                                                .readdata
		.player1Score0_s1_writedata                                            (mm_interconnect_0_player1score0_s1_writedata),                //                                                                .writedata
		.player1Score0_s1_chipselect                                           (mm_interconnect_0_player1score0_s1_chipselect),               //                                                                .chipselect
		.player1Score1_s1_address                                              (mm_interconnect_0_player1score1_s1_address),                  //                                                player1Score1_s1.address
		.player1Score1_s1_write                                                (mm_interconnect_0_player1score1_s1_write),                    //                                                                .write
		.player1Score1_s1_readdata                                             (mm_interconnect_0_player1score1_s1_readdata),                 //                                                                .readdata
		.player1Score1_s1_writedata                                            (mm_interconnect_0_player1score1_s1_writedata),                //                                                                .writedata
		.player1Score1_s1_chipselect                                           (mm_interconnect_0_player1score1_s1_chipselect),               //                                                                .chipselect
		.player2Score0_s1_address                                              (mm_interconnect_0_player2score0_s1_address),                  //                                                player2Score0_s1.address
		.player2Score0_s1_write                                                (mm_interconnect_0_player2score0_s1_write),                    //                                                                .write
		.player2Score0_s1_readdata                                             (mm_interconnect_0_player2score0_s1_readdata),                 //                                                                .readdata
		.player2Score0_s1_writedata                                            (mm_interconnect_0_player2score0_s1_writedata),                //                                                                .writedata
		.player2Score0_s1_chipselect                                           (mm_interconnect_0_player2score0_s1_chipselect),               //                                                                .chipselect
		.player2Score1_s1_address                                              (mm_interconnect_0_player2score1_s1_address),                  //                                                player2Score1_s1.address
		.player2Score1_s1_write                                                (mm_interconnect_0_player2score1_s1_write),                    //                                                                .write
		.player2Score1_s1_readdata                                             (mm_interconnect_0_player2score1_s1_readdata),                 //                                                                .readdata
		.player2Score1_s1_writedata                                            (mm_interconnect_0_player2score1_s1_writedata),                //                                                                .writedata
		.player2Score1_s1_chipselect                                           (mm_interconnect_0_player2score1_s1_chipselect),               //                                                                .chipselect
		.sdram_s1_address                                                      (mm_interconnect_0_sdram_s1_address),                          //                                                        sdram_s1.address
		.sdram_s1_write                                                        (mm_interconnect_0_sdram_s1_write),                            //                                                                .write
		.sdram_s1_read                                                         (mm_interconnect_0_sdram_s1_read),                             //                                                                .read
		.sdram_s1_readdata                                                     (mm_interconnect_0_sdram_s1_readdata),                         //                                                                .readdata
		.sdram_s1_writedata                                                    (mm_interconnect_0_sdram_s1_writedata),                        //                                                                .writedata
		.sdram_s1_byteenable                                                   (mm_interconnect_0_sdram_s1_byteenable),                       //                                                                .byteenable
		.sdram_s1_readdatavalid                                                (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                                                .readdatavalid
		.sdram_s1_waitrequest                                                  (mm_interconnect_0_sdram_s1_waitrequest),                      //                                                                .waitrequest
		.sdram_s1_chipselect                                                   (mm_interconnect_0_sdram_s1_chipselect),                       //                                                                .chipselect
		.sdram_pll_audio_pll_pll_slave_address                                 (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_address),     //                                   sdram_pll_audio_pll_pll_slave.address
		.sdram_pll_audio_pll_pll_slave_write                                   (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_write),       //                                                                .write
		.sdram_pll_audio_pll_pll_slave_read                                    (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_read),        //                                                                .read
		.sdram_pll_audio_pll_pll_slave_readdata                                (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_readdata),    //                                                                .readdata
		.sdram_pll_audio_pll_pll_slave_writedata                               (mm_interconnect_0_sdram_pll_audio_pll_pll_slave_writedata),   //                                                                .writedata
		.sysid_qsys_0_control_slave_address                                    (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //                                      sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                   (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                                                .readdata
		.timer_0_s1_address                                                    (mm_interconnect_0_timer_0_s1_address),                        //                                                      timer_0_s1.address
		.timer_0_s1_write                                                      (mm_interconnect_0_timer_0_s1_write),                          //                                                                .write
		.timer_0_s1_readdata                                                   (mm_interconnect_0_timer_0_s1_readdata),                       //                                                                .readdata
		.timer_0_s1_writedata                                                  (mm_interconnect_0_timer_0_s1_writedata),                      //                                                                .writedata
		.timer_0_s1_chipselect                                                 (mm_interconnect_0_timer_0_s1_chipselect),                     //                                                                .chipselect
		.timeScreen0_s1_address                                                (mm_interconnect_0_timescreen0_s1_address),                    //                                                  timeScreen0_s1.address
		.timeScreen0_s1_write                                                  (mm_interconnect_0_timescreen0_s1_write),                      //                                                                .write
		.timeScreen0_s1_readdata                                               (mm_interconnect_0_timescreen0_s1_readdata),                   //                                                                .readdata
		.timeScreen0_s1_writedata                                              (mm_interconnect_0_timescreen0_s1_writedata),                  //                                                                .writedata
		.timeScreen0_s1_chipselect                                             (mm_interconnect_0_timescreen0_s1_chipselect),                 //                                                                .chipselect
		.timeScreen1_s1_address                                                (mm_interconnect_0_timescreen1_s1_address),                    //                                                  timeScreen1_s1.address
		.timeScreen1_s1_write                                                  (mm_interconnect_0_timescreen1_s1_write),                      //                                                                .write
		.timeScreen1_s1_readdata                                               (mm_interconnect_0_timescreen1_s1_readdata),                   //                                                                .readdata
		.timeScreen1_s1_writedata                                              (mm_interconnect_0_timescreen1_s1_writedata),                  //                                                                .writedata
		.timeScreen1_s1_chipselect                                             (mm_interconnect_0_timescreen1_s1_chipselect),                 //                                                                .chipselect
		.timeScreen2_s1_address                                                (mm_interconnect_0_timescreen2_s1_address),                    //                                                  timeScreen2_s1.address
		.timeScreen2_s1_write                                                  (mm_interconnect_0_timescreen2_s1_write),                      //                                                                .write
		.timeScreen2_s1_readdata                                               (mm_interconnect_0_timescreen2_s1_readdata),                   //                                                                .readdata
		.timeScreen2_s1_writedata                                              (mm_interconnect_0_timescreen2_s1_writedata),                  //                                                                .writedata
		.timeScreen2_s1_chipselect                                             (mm_interconnect_0_timescreen2_s1_chipselect)                  //                                                                .chipselect
	);

	Bomberman_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_qsys_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_audio_pll_c0_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
